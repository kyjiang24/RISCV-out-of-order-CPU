`ifndef MACROS_SVH  // header guard to prevent multiple include error
`define MACROS_SVH

`define BENCHMARK "test_sb_type"
`define SIM_CYCLES 800                   // change number of cycles to run simulation for
`define TESTING_NON_SYNTH               // comment out to disable automated testing

// define commonly used constants
`define example 2'b00

`endif  // MACROS_SVH
